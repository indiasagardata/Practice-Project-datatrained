# Practice-Project-datatrained

https://indiasagardata.github.io/Practice-Project-datatrained/ tap here to quick preview my work
